`include "ternary_logic.v"

module testbench();

  reg x = 0;
  reg y = 0;
  reg w = 0;
  reg v = 0;
  wire z;
  wire and_out;
  wire or_out;
//  wire [1:0] c; // Изменили тип порта c на wire
  wire and_result;
  wire nand_result;
  wire not_out;
  wire clos_out;
  wire not_v_out;
  wire not_y_out;
  wire s;
  not_gate not_v(v, not_v_out);
  not_gate not_y(y, not_y_out);
  and_4_gate clos_h(x, not_y_out, w, not_v_out, clos_out);

  and_4_gate nand_xy(x, y, w, v, z);
  or_gate or_xy(x, y, or_out);
  and_gate and_xy(x, y, and_out);
  not_gate not_x(x, not_out);
  initial begin
    $display("and_4_gate: ");
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 0; y = 0; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 0; y = 0; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 0; y = 0; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 0; y = 1; w = 0; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 0; y = 1; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 0; y = 1; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 0; y = 1; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 0; w = 0; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 0; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 0; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 0; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 1; w = 0; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 1; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 1; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    #5 x = 1; y = 1; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, z);
    $display("or_gate: ");
    #5 x = 0; y = 0;
    $display("x = %b, y = %b,z = %b", x, y, or_out);
    #5 x = 0; y = 1;
    $display("x = %b, y = %b,z = %b", x, y, or_out);
    #5 x = 1; y = 0;
    $display("x = %b, y = %b,z = %b", x, y, or_out);
    #5 x = 1; y = 1;
    $display("x = %b, y = %b,z = %b", x, y, or_out);
    $display("and_gate: ");
    #5 x = 0; y = 0;
    $display("x = %b, y = %b,z = %b", x, y, and_out);
    #5 x = 0; y = 1;
    $display("x = %b, y = %b,z = %b", x, y, and_out);
    #5 x = 1; y = 0;
    $display("x = %b, y = %b,z = %b", x, y, and_out);
    #5 x = 1; y = 1;
    $display("x = %b, y = %b,z = %b", x, y, and_out);
    $display("not_gate: ");
    #5 x = 0; 
    $display("x = %b,z = %b", x, not_out);
    #5 x = 1; 
    $display("x = %b,z = %b", x, not_out);
    $display("and_4_gate_clos: ");
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 0; y = 0; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 0; y = 0; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 0; y = 0; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 0; y = 1; w = 0; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 0; y = 1; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 0; y = 1; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 0; y = 1; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 0; w = 0; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 0; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 0; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 0; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 1; w = 0; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 1; w = 0; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 1; w = 1; v = 0;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);
    #5 x = 1; y = 1; w = 1; v = 1;  
    $display("x = %b, y = %b, w = %b, v = %b, z = %b", x, y, w, v, clos_out);

  end
endmodule